library verilog;
use verilog.vl_types.all;
entity Imem_vlg_vec_tst is
end Imem_vlg_vec_tst;
