library verilog;
use verilog.vl_types.all;
entity MEMORY_vlg_vec_tst is
end MEMORY_vlg_vec_tst;
