library verilog;
use verilog.vl_types.all;
entity EXECUTE_vlg_vec_tst is
end EXECUTE_vlg_vec_tst;
