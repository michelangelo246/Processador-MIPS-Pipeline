library verilog;
use verilog.vl_types.all;
entity DECODE_vlg_vec_tst is
end DECODE_vlg_vec_tst;
