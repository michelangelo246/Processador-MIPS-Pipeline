library verilog;
use verilog.vl_types.all;
entity FETCH_vlg_vec_tst is
end FETCH_vlg_vec_tst;
