library verilog;
use verilog.vl_types.all;
entity ULA_vlg_vec_tst is
end ULA_vlg_vec_tst;
