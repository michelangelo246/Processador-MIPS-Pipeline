library verilog;
use verilog.vl_types.all;
entity MemI_vlg_vec_tst is
end MemI_vlg_vec_tst;
