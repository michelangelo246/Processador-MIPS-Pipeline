library verilog;
use verilog.vl_types.all;
entity ControleULA_vlg_vec_tst is
end ControleULA_vlg_vec_tst;
